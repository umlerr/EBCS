library verilog;
use verilog.vl_types.all;
entity Pract2_Misha_vlg_sample_tst is
    port(
        x_1             : in     vl_logic;
        x_2             : in     vl_logic;
        x_3             : in     vl_logic;
        x_4             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Pract2_Misha_vlg_sample_tst;
