library verilog;
use verilog.vl_types.all;
entity music_project_vlg_vec_tst is
end music_project_vlg_vec_tst;
