library verilog;
use verilog.vl_types.all;
entity lab1_vlg_check_tst is
    port(
        y_and           : in     vl_logic;
        y_or            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab1_vlg_check_tst;
