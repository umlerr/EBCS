library verilog;
use verilog.vl_types.all;
entity Pract2_Misha is
    port(
        y               : out    vl_logic;
        x_1             : in     vl_logic;
        x_2             : in     vl_logic;
        x_3             : in     vl_logic;
        x_4             : in     vl_logic;
        \1Y\            : out    vl_logic;
        \2Y\            : out    vl_logic
    );
end Pract2_Misha;
