library verilog;
use verilog.vl_types.all;
entity tmp_vlg_check_tst is
    port(
        D0              : in     vl_logic;
        D00             : in     vl_logic;
        D1              : in     vl_logic;
        D01             : in     vl_logic;
        D2              : in     vl_logic;
        D02             : in     vl_logic;
        D3              : in     vl_logic;
        D03             : in     vl_logic;
        D4              : in     vl_logic;
        D04             : in     vl_logic;
        D5              : in     vl_logic;
        D05             : in     vl_logic;
        D6              : in     vl_logic;
        D06             : in     vl_logic;
        DP              : in     vl_logic;
        y0              : in     vl_logic;
        y1              : in     vl_logic;
        y2              : in     vl_logic;
        y3              : in     vl_logic;
        y4              : in     vl_logic;
        y5              : in     vl_logic;
        y6              : in     vl_logic;
        y7              : in     vl_logic;
        y8              : in     vl_logic;
        y9              : in     vl_logic;
        y10             : in     vl_logic;
        y11             : in     vl_logic;
        y12             : in     vl_logic;
        y13             : in     vl_logic;
        y14             : in     vl_logic;
        y15             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end tmp_vlg_check_tst;
