library verilog;
use verilog.vl_types.all;
entity tmp is
    port(
        D0              : out    vl_logic;
        y1              : out    vl_logic;
        x               : in     vl_logic_vector(3 downto 0);
        y11             : out    vl_logic;
        y4              : out    vl_logic;
        y14             : out    vl_logic;
        D1              : out    vl_logic;
        y5              : out    vl_logic;
        y6              : out    vl_logic;
        y15             : out    vl_logic;
        D2              : out    vl_logic;
        y12             : out    vl_logic;
        y2              : out    vl_logic;
        D3              : out    vl_logic;
        y7              : out    vl_logic;
        D4              : out    vl_logic;
        y13             : out    vl_logic;
        y3              : out    vl_logic;
        y9              : out    vl_logic;
        D5              : out    vl_logic;
        D6              : out    vl_logic;
        y0              : out    vl_logic;
        y10             : out    vl_logic;
        DP              : out    vl_logic;
        D00             : out    vl_logic;
        D01             : out    vl_logic;
        D02             : out    vl_logic;
        D03             : out    vl_logic;
        D04             : out    vl_logic;
        D05             : out    vl_logic;
        D06             : out    vl_logic;
        y8              : out    vl_logic
    );
end tmp;
