library verilog;
use verilog.vl_types.all;
entity RS_trigger_vlg_vec_tst is
end RS_trigger_vlg_vec_tst;
