library verilog;
use verilog.vl_types.all;
entity Lab7_3 is
    port(
        D               : out    vl_logic_vector(3 downto 0);
        C               : in     vl_logic
    );
end Lab7_3;
