library verilog;
use verilog.vl_types.all;
entity lab2_1_vlg_check_tst is
    port(
        dec_out         : in     vl_logic;
        lab1_out        : in     vl_logic;
        mux_out         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab2_1_vlg_check_tst;
