library verilog;
use verilog.vl_types.all;
entity Coursework_mux_vlg_vec_tst is
end Coursework_mux_vlg_vec_tst;
