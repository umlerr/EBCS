library verilog;
use verilog.vl_types.all;
entity Coursework_vlg_vec_tst is
end Coursework_vlg_vec_tst;
