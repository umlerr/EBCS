library verilog;
use verilog.vl_types.all;
entity kurs_vlg_sample_tst is
    port(
        C               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end kurs_vlg_sample_tst;
