library verilog;
use verilog.vl_types.all;
entity Lab5_2_vlg_vec_tst is
end Lab5_2_vlg_vec_tst;
