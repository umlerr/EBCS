library verilog;
use verilog.vl_types.all;
entity lab2_1_vlg_vec_tst is
end lab2_1_vlg_vec_tst;
