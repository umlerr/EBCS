library verilog;
use verilog.vl_types.all;
entity Lab6_1_vlg_vec_tst is
end Lab6_1_vlg_vec_tst;
