library verilog;
use verilog.vl_types.all;
entity Lab7_1_vlg_vec_tst is
end Lab7_1_vlg_vec_tst;
