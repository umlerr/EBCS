library verilog;
use verilog.vl_types.all;
entity Pract2_vlg_vec_tst is
end Pract2_vlg_vec_tst;
