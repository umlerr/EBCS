library verilog;
use verilog.vl_types.all;
entity kurs_vlg_vec_tst is
end kurs_vlg_vec_tst;
