library verilog;
use verilog.vl_types.all;
entity tmp_vlg_vec_tst is
end tmp_vlg_vec_tst;
