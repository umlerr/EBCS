library verilog;
use verilog.vl_types.all;
entity Pract2 is
    port(
        \out\           : out    vl_logic;
        x               : in     vl_logic_vector(3 downto 0)
    );
end Pract2;
