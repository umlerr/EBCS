library verilog;
use verilog.vl_types.all;
entity Lab6_2_vlg_vec_tst is
end Lab6_2_vlg_vec_tst;
