library verilog;
use verilog.vl_types.all;
entity JK_trigger_vlg_vec_tst is
end JK_trigger_vlg_vec_tst;
