library verilog;
use verilog.vl_types.all;
entity Lab7_2_vlg_sample_tst is
    port(
        C               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Lab7_2_vlg_sample_tst;
